module sample(
  input x,
  input y,
  output sum
)
assign sum = x + y;
endmodule
